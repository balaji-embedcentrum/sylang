circuit ControlSignalCircuit
  name "Control Signal Output Circuit"  
  description "Electronics circuit for digital control outputs including backup enable and actuator type selection with safety interlocks and diagnostics"
  owner "Electronics Team"
  tags "control", "digital-output", "backup", "selection"
  safetylevel ASIL-D
  partof ActuatorManagementUnit
  
  implements BackupActivationController
  
  interfaces
    Backup_Enable "3.3V CMOS digital output"
    Actuator_Type_Select "4-bit digital output selection" 