circuit CommunicationCircuit
  name "Automation Communication Circuit"
  description "Electronics circuit for automation communication interfaces, data exchange, and system coordination signals"
  owner "Electronics Team"
  tags "communication", "coordination", "data-exchange", "interfaces"
  safetylevel ASIL-B
  partof AutomationCoordinationUnit
  
  interfaces
    System_Communication_Bus "System-wide communication bus interface"
    Coordination_Data_Exchange "Component coordination data interface"
    Status_Reporting_Interface "Automation status reporting interface" 