electronicscircuit EthernetInterfaceCircuit
  name "Ethernet Interface Circuit"
  description "Electronics circuit providing Ethernet PHY functionality, frame processing, and TSN hardware support"
  owner "Electronics Team"
  tags "Ethernet-interface", "PHY", "frame-processing", "TSN-hardware"
  safetylevel ASIL-B
  partof StandardsComplianceUnit
  implements EthernetFrameProcessor, TSNConfigurationEngine
  interfaces
    input ethernet_signals "Ethernet differential signals and network data streams"
    input ethernet_control_signals "Ethernet PHY control signals and configuration commands"
    output ethernet_phy "Ethernet PHY functionality and signal processing"
    output ethernet_frame_processor "Hardware Ethernet frame processing and packet handling"
    output tsn_hardware "Time-Sensitive Networking hardware support and real-time control"
