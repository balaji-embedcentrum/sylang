circuit CurrentSensingCircuit
  name "Current Sensing Circuit"
  description "Electronics circuit for motor current sensing, measurement conditioning, and overcurrent protection"
  owner "Electronics Team"
  tags "current", "sensing", "measurement", "protection"
  safetylevel ASIL-D
  partof MotorControlUnit
  
  implements CurrentSensingProcessor
  
  interfaces
    Current_Sensor_Input "Current sensor measurement inputs"
    Current_Measurement_Output "Conditioned current measurements"
    Overcurrent_Protection "Overcurrent protection signals" 