circuit PowerDistributionCircuit
  name "Power Distribution Circuit"
  description "Electronics circuit for power distribution, load switching, and power allocation management"
  owner "Electronics Team"
  tags "power", "distribution", "switching", "allocation"
  safetylevel ASIL-D
  partof PowerManagementUnit
  
  implements PowerDistributionController
  
  interfaces
    Power_Input "Main power input"
    Distributed_Outputs "Multiple power distribution outputs"
    Load_Control "Load switching control signals" 