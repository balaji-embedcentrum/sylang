circuit AutomationControlCircuit
  name "Automation Control Circuit"
  description "Electronics circuit for automation control signals, state machine processing, and arbitration control interfaces"
  owner "Electronics Team"
  tags "automation", "control", "state-machine", "arbitration"
  safetylevel ASIL-B
  partof AutomationCoordinationUnit
  
  implements StateTransitionController, ActivationSequencer, RequestPriorityManager
  
  interfaces
    Automation_Control_Input "Automation control signal inputs"
    State_Control_Output "State machine control outputs"
    Priority_Control_Output "Request priority control signals" 