circuit PowerElectronicsCircuit
  name "Power Electronics Circuit"
  description "Electronics circuit for motor power electronics, inverter control, and high-voltage power switching"
  owner "Electronics Team"
  tags "power", "electronics", "inverter", "switching"
  safetylevel ASIL-D
  partof MotorControlUnit
  
  interfaces
    High_Voltage_Input "High voltage power input"
    Inverter_Control "Inverter switching control"
    Power_Protection "Power electronics protection" 